`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2026/01/19 02:08:35
// Design Name: 
// Module Name: top
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module top(
    input CLK, // ������ʱ�ӣ�ϵͳʱ��
    input RST, // �͵�ƽ��Ч��λ
    // MP3����JC
    input DREQ,      // VS1003 ���������ź�
    output XDCS, // ����Ƭѡ
    output XCS,  // ����Ƭѡ
    output RSET, 
    output SI,   // ��������
    output SCLK,  // VS1003 ʱ��
    // ����
    input BTNC,
    input BTNU,
    input BTND,
    input BTNL,
    input BTNR,
    // ��������ֱ��ѡ�����
    input [15:0] SW,
    // 7 �������
    output [6: 0] SEG,
    output [7: 0] SHIFT,
    output DOT,
    // OLED �ӿڣ���JB
    output DIN,
    output OLED_CLK,
    output CS,
    output DC,
    output RES,
    // ������ʾ LED
    output [15: 0] led
);
    wire [15:0] vol_code_bus;  // �������ɰ���ģ��������
    wire [2:0] song_idx_bus;// ��ǰ����������Ŀǰ���8��
    reg [15:0] elapsed_secs;// ʱ����� (��)
    integer clk_ticks_count; // ��ʱ�Ӽ����������뼶�ۼ�
    wire mp3_rst_sync; // ���� MP3 �ĸ�λ/��ʾ��λ�ź�
     // 7 ���������ʾ
       Display7 u_seg7_display(
           .CLK(CLK),
           .DATA(elapsed_secs),
           .VOL(vol_code_bus),
           .CURRENT(song_idx_bus),
           .SEG(SEG),
           .SHIFT(SHIFT),
           .DOT(DOT)
       );
    // ��������
    btn_control u_button_ctrl(
        .CLK(CLK),
        .RST(RST),
        .BTNC(BTNC),
        .BTNU(BTNU),
        .BTND(BTND),
        .BTNL(BTNL),
        .BTNR(BTNR),
        .SW(SW),
        .vol(vol_code_bus),
        .CURRENT(song_idx_bus)
    );
    // OLED ģ��
    oled u_oled_display(
        .CLK(CLK), 
        .RST(RST),
        .current(song_idx_bus),
        .DIN(DIN),
        .OLED_CLK(OLED_CLK), 
        .CS(CS),
        .DC(DC),
        .RES(RES)
    );
    // MP3 ģ��
    MP3 u_mp3_player(
        .CLK(CLK), 
        .RST(RST), 
        .DREQ(DREQ),
        .vol(vol_code_bus),
        .current(song_idx_bus),
        .XDCS(XDCS), 
        .XCS(XCS), 
        .RSET(RSET), 
        .SI(SI),
        .SCLK(SCLK),
        .MP3_RST(mp3_rst_sync),
        .led(led)
    );
    //����������ģ��
    always @ (posedge CLK) begin
        if(!RST) begin
            elapsed_secs <= 16'd0;
            clk_ticks_count <= 0;
        end else if((clk_ticks_count+1)==100000000) begin
            clk_ticks_count <= 0;
            elapsed_secs <= elapsed_secs + 1;
        end else begin
            clk_ticks_count <= clk_ticks_count + 1;
        end
    end
endmodule
